CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 230 30 400 10
176 80 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 40 334 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-32 -6 -18 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44797.6 0
0
13 Logic Switch~
5 40 407 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-32 2 -18 10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44797.6 0
0
13 Logic Switch~
5 83 221 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-36 1 -22 9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
44797.6 0
0
13 Logic Switch~
5 100 152 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-43 -2 -29 6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
44797.6 0
0
13 Logic Switch~
5 100 95 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-40 -3 -26 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
44797.6 0
0
14 Logic Display~
6 253 406 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
44797.6 0
0
14 Logic Display~
6 238 317 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
44797.6 0
0
9 Inverter~
13 92 379 0 2 22
0 4 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
7361 0 0
2
44797.6 0
0
5 4081~
219 173 416 0 3 22
0 4 5 2
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
4747 0 0
2
44797.6 0
0
5 4081~
219 163 336 0 3 22
0 6 5 3
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
972 0 0
2
44797.6 0
0
9 Inverter~
13 133 215 0 2 22
0 8 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3472 0 0
2
44797.6 0
0
14 Logic Display~
6 326 127 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
44797.6 0
0
5 4071~
219 245 133 0 3 22
0 11 10 7
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3536 0 0
2
44797.6 0
0
5 4081~
219 162 162 0 3 22
0 12 9 10
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
4597 0 0
2
44797.6 0
0
5 4081~
219 162 108 0 3 22
0 13 8 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3835 0 0
2
44797.6 0
0
15
3 1 2 0 0 4224 0 9 6 0 0 4
194 416
235 416
235 424
253 424
3 1 3 0 0 8320 0 10 7 0 0 3
184 336
184 335
238 335
0 1 4 0 0 4096 0 0 8 4 0 3
61 407
61 379
77 379
1 1 4 0 0 4224 0 2 9 0 0 2
52 407
149 407
1 2 5 0 0 4096 0 1 9 0 0 5
52 334
52 392
99 392
99 425
149 425
2 1 6 0 0 4224 0 8 10 0 0 3
113 379
113 327
139 327
1 2 5 0 0 4224 0 1 10 0 0 4
52 334
116 334
116 345
139 345
3 1 7 0 0 4224 0 13 12 0 0 4
278 133
312 133
312 145
326 145
0 2 8 0 0 4224 0 0 15 10 0 3
111 215
111 117
138 117
1 1 8 0 0 0 0 3 11 0 0 4
95 221
111 221
111 215
118 215
2 2 9 0 0 4224 0 11 14 0 0 5
154 215
154 183
129 183
129 171
138 171
3 2 10 0 0 4224 0 14 13 0 0 4
183 162
215 162
215 142
232 142
3 1 11 0 0 4224 0 15 13 0 0 4
183 108
214 108
214 124
232 124
1 1 12 0 0 8320 0 4 14 0 0 3
112 152
112 153
138 153
1 1 13 0 0 4224 0 5 15 0 0 4
112 95
130 95
130 99
138 99
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
41 267 152 291
44 269 148 285
13 Demultiplexor
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
83 58 178 82
86 60 174 76
11 multiplexor
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
