CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
36
5 4071~
219 739 241 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
7361 0 0
2
44795.7 0
0
5 4071~
219 818 287 0 3 22
0 25 24 23
0
0 0 96 0
4 4071
-7 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
4747 0 0
2
44795.7 5
0
9 Inverter~
13 912 288 0 2 22
0 23 22
0
0 0 96 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
972 0 0
2
44795.7 4
0
14 Logic Display~
6 957 269 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
44795.7 3
0
13 Logic Switch~
5 669 217 0 1 11
0 27
0
0 0 21344 0
2 0V
-5 -16 9 -8
1 A
-30 -4 -23 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9998 0 0
2
44795.7 2
0
13 Logic Switch~
5 668 269 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 B
-31 -5 -24 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3536 0 0
2
44795.7 1
0
13 Logic Switch~
5 669 319 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-5 -16 9 -8
1 C
-31 -4 -24 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4597 0 0
2
44795.7 0
0
13 Logic Switch~
5 158 951 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-27 -3 -20 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3835 0 0
2
44795.7 4
0
13 Logic Switch~
5 159 1059 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-28 -1 -21 7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3670 0 0
2
44795.7 3
0
13 Logic Switch~
5 159 1112 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-26 -3 -19 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5616 0 0
2
44795.7 2
0
13 Logic Switch~
5 157 1158 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-30 -4 -23 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9323 0 0
2
44795.7 1
0
13 Logic Switch~
5 153 1207 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 E
-29 2 -22 10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
317 0 0
2
44795.7 0
0
13 Logic Switch~
5 131 724 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 E
-31 1 -24 9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3108 0 0
2
44795.6 0
0
13 Logic Switch~
5 139 672 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-30 -4 -23 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4299 0 0
2
44795.6 0
0
13 Logic Switch~
5 144 626 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-26 -3 -19 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9672 0 0
2
44795.6 0
0
13 Logic Switch~
5 143 578 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-28 -1 -21 7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7876 0 0
2
44795.6 0
0
13 Logic Switch~
5 142 495 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-27 -3 -20 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6369 0 0
2
44795.6 0
0
13 Logic Switch~
5 106 317 0 1 11
0 24
0
0 0 21360 0
2 0V
-5 -16 9 -8
1 C
-31 -4 -24 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9172 0 0
2
44795.6 0
0
13 Logic Switch~
5 105 267 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-31 -5 -24 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7100 0 0
2
44795.6 0
0
13 Logic Switch~
5 106 215 0 1 11
0 27
0
0 0 21360 0
2 0V
-5 -16 9 -8
1 A
-30 -4 -23 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3820 0 0
2
44795.6 0
0
5 4071~
219 516 1069 0 3 22
0 6 5 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
7678 0 0
2
44795.7 0
0
5 4071~
219 261 1008 0 3 22
0 11 10 8
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
961 0 0
2
44795.7 10
0
5 4081~
219 361 1062 0 3 22
0 8 9 7
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3178 0 0
2
44795.7 9
0
9 Inverter~
13 438 1061 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3409 0 0
2
44795.7 8
0
5 4081~
219 627 1120 0 3 22
0 2 4 3
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3951 0 0
2
44795.7 6
0
14 Logic Display~
6 686 1102 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8885 0 0
2
44795.7 5
0
14 Logic Display~
6 670 621 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3780 0 0
2
44795.6 0
0
5 4081~
219 611 639 0 3 22
0 14 13 12
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
9265 0 0
2
44795.6 0
0
6 74266~
219 501 588 0 3 22
0 16 15 14
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9442 0 0
2
44795.6 0
0
9 Inverter~
13 422 580 0 2 22
0 17 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
9424 0 0
2
44795.6 0
0
5 4081~
219 345 581 0 3 22
0 18 19 17
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9968 0 0
2
44795.6 0
0
5 4071~
219 245 527 0 3 22
0 21 20 18
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9281 0 0
2
44795.6 0
0
14 Logic Display~
6 394 267 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8464 0 0
2
44795.6 0
0
9 Inverter~
13 349 286 0 2 22
0 23 22
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
7168 0 0
2
44795.6 0
0
5 4071~
219 255 285 0 3 22
0 25 24 23
0
0 0 112 0
4 4071
-7 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3171 0 0
2
44795.6 0
0
5 4081~
219 188 239 0 3 22
0 27 26 25
0
0 0 112 0
4 4081
-7 -24 21 -16
0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
4139 0 0
2
44795.6 0
0
32
2 1 22 0 0 16 0 3 4 0 0 3
933 288
933 287
957 287
3 1 23 0 0 16 0 2 3 0 0 3
851 287
851 288
897 288
1 2 24 0 0 16 0 7 2 0 0 4
681 319
785 319
785 296
805 296
3 1 25 0 0 16 0 1 2 0 0 3
772 241
805 241
805 278
1 2 26 0 0 16 0 6 1 0 0 4
680 269
727 269
727 250
726 250
1 1 27 0 0 16 0 5 1 0 0 4
681 217
727 217
727 232
726 232
3 1 2 0 0 4224 0 21 25 0 0 3
549 1069
603 1069
603 1111
3 1 3 0 0 4224 0 25 26 0 0 2
648 1120
686 1120
1 2 4 0 0 4224 0 12 25 0 0 3
165 1207
603 1207
603 1129
1 2 5 0 0 4224 0 11 21 0 0 4
169 1158
501 1158
501 1078
503 1078
2 1 6 0 0 8320 0 24 21 0 0 3
459 1061
459 1060
503 1060
3 1 7 0 0 8320 0 23 24 0 0 3
382 1062
382 1061
423 1061
3 1 8 0 0 8320 0 22 23 0 0 3
294 1008
337 1008
337 1053
1 2 9 0 0 4224 0 10 23 0 0 3
171 1112
337 1112
337 1071
1 2 10 0 0 4224 0 9 22 0 0 3
171 1059
248 1059
248 1017
1 1 11 0 0 4224 0 8 22 0 0 3
170 951
248 951
248 999
3 1 12 0 0 4224 0 28 27 0 0 2
632 639
670 639
1 2 13 0 0 4224 0 13 28 0 0 3
143 724
587 724
587 648
3 1 14 0 0 4224 0 29 28 0 0 3
540 588
587 588
587 630
1 2 15 0 0 4224 0 14 29 0 0 3
151 672
485 672
485 597
2 1 16 0 0 8320 0 30 29 0 0 3
443 580
443 579
485 579
3 1 17 0 0 8320 0 31 30 0 0 3
366 581
366 580
407 580
3 1 18 0 0 8320 0 32 31 0 0 3
278 527
321 527
321 572
1 2 19 0 0 4224 0 15 31 0 0 3
156 626
321 626
321 590
1 2 20 0 0 4224 0 16 32 0 0 3
155 578
232 578
232 536
1 1 21 0 0 4224 0 17 32 0 0 3
154 495
232 495
232 518
2 1 22 0 0 8320 0 34 33 0 0 3
370 286
370 285
394 285
3 1 23 0 0 8320 0 35 34 0 0 3
288 285
288 286
334 286
1 2 24 0 0 4224 0 18 35 0 0 4
118 317
222 317
222 294
242 294
3 1 25 0 0 8320 0 36 35 0 0 3
209 239
242 239
242 276
1 2 26 0 0 4224 0 19 36 0 0 3
117 267
164 267
164 248
1 1 27 0 0 4224 0 20 36 0 0 3
118 215
164 215
164 230
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
