CircuitMaker Text
5.6
Probes: 1
v2[p]
Transient Analysis
0 255 87 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 110 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 1532 488
9437202 0
0
6 Title:
5 Name:
0
0
0
8
2 +V
167 256 68 0 1 3
0 4
0
0 0 54384 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
5 OUPUT
-16 -14 19 -6
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5130 0 0
2
44803.8 0
0
7 Ground~
168 317 575 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
391 0 0
2
44803.8 0
0
2 +V
167 401 122 0 1 3
0 3
0
0 0 54256 0
2 9V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3124 0 0
2
44803.8 0
0
10 Capacitor~
219 439 513 0 2 5
0 2 7
0
0 0 848 90
3 1nF
11 0 32 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
3421 0 0
2
44803.8 0
0
10 555 Timer~
219 379 335 0 8 17
0 2 6 4 3 7 6 5 3
0
0 0 4944 0
3 555
-11 -36 10 -28
2 U1
-7 -46 7 -38
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 0 0 0 0 0
1 U
8157 0 0
2
44803.8 0
0
10 Capacitor~
219 115 529 0 2 5
0 2 6
0
0 0 848 90
4 47uF
12 0 40 8
2 C1
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
5572 0 0
2
44803.8 0
0
9 Resistor~
219 115 424 0 2 5
0 6 5
0
0 0 880 90
3 50k
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8901 0 0
2
44803.8 0
0
9 Resistor~
219 114 156 0 4 5
0 5 3 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7361 0 0
2
44803.8 0
0
13
1 1 2 0 0 4224 0 2 5 0 0 3
317 569
317 326
347 326
1 1 2 0 0 0 0 2 4 0 0 3
317 569
439 569
439 522
1 1 2 0 0 0 0 6 2 0 0 3
115 538
115 569
317 569
0 8 3 0 0 4096 0 0 5 7 0 4
401 138
401 288
411 288
411 326
1 3 4 0 0 4224 0 1 5 0 0 3
256 77
256 344
347 344
0 4 3 0 0 4096 0 0 5 7 0 3
166 138
166 353
347 353
2 1 3 0 0 4224 0 8 3 0 0 3
114 138
401 138
401 131
0 7 5 0 0 12416 0 0 5 13 0 6
115 367
177 367
177 393
457 393
457 335
411 335
0 2 6 0 0 12288 0 0 5 10 0 4
218 419
241 419
241 335
347 335
0 6 6 0 0 12416 0 0 5 12 0 6
115 461
218 461
218 374
451 374
451 344
411 344
5 2 7 0 0 8320 0 5 4 0 0 3
411 353
439 353
439 504
1 2 6 0 0 0 0 7 6 0 0 2
115 442
115 520
1 2 5 0 0 0 0 8 7 0 0 3
114 174
115 174
115 406
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
