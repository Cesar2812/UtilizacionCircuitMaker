CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 430 30 400 10
176 80 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
32
13 Logic Switch~
5 42 602 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 E
-30 -5 -23 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44795.7 0
0
13 Logic Switch~
5 41 564 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 D
-32 -3 -25 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44795.7 0
0
13 Logic Switch~
5 42 530 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-29 -2 -22 6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44795.7 0
0
13 Logic Switch~
5 42 497 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-27 -3 -20 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
44795.7 0
0
13 Logic Switch~
5 42 467 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-29 -3 -22 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
44795.7 0
0
13 Logic Switch~
5 99 419 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-28 -4 -21 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5572 0 0
2
44795.6 0
0
13 Logic Switch~
5 97 372 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-26 -3 -19 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
44795.6 0
0
13 Logic Switch~
5 95 324 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-26 -5 -19 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
44795.6 0
0
13 Logic Switch~
5 95 284 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-28 -4 -21 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4747 0 0
2
44795.6 0
0
13 Logic Switch~
5 94 234 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-25 -4 -18 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
972 0 0
2
44795.6 0
0
13 Logic Switch~
5 94 186 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-27 -4 -20 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3472 0 0
2
44795.6 0
0
13 Logic Switch~
5 87 128 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-9 10 5 18
1 C
-27 -4 -20 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
5.90044e-315 0
0
13 Logic Switch~
5 87 56 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-23 -4 -16 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90044e-315 0
0
13 Logic Switch~
5 88 91 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
1 B
-25 -6 -18 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
5.90044e-315 0
0
14 Logic Display~
6 458 550 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
44795.7 0
0
5 4081~
219 393 563 0 3 22
0 3 4 2
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndD
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3670 0 0
2
44795.7 0
0
5 4030~
219 320 534 0 3 22
0 5 6 3
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
5616 0 0
2
44795.7 0
0
9 Inverter~
13 248 517 0 2 22
0 7 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
9323 0 0
2
44795.7 0
0
5 4081~
219 173 517 0 3 22
0 8 9 7
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndC
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
317 0 0
2
44795.7 0
0
5 4071~
219 101 483 0 3 22
0 11 10 8
0
0 0 624 0
4 4071
-7 -24 21 -16
3 OrD
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3108 0 0
2
44795.7 0
0
14 Logic Display~
6 327 361 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
44795.7 0
0
5 4073~
219 171 398 0 4 22
0 17 16 15 13
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
9672 0 0
2
44795.7 0
0
5 4023~
219 155 344 0 4 22
0 17 16 15 14
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 4 0
1 U
7876 0 0
2
44795.7 0
0
5 4071~
219 264 374 0 3 22
0 14 13 12
0
0 0 624 0
4 4071
-7 -24 21 -16
3 OrC
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
6369 0 0
2
44795.7 0
0
14 Logic Display~
6 351 231 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9172 0 0
2
44795.6 0
0
9 Inverter~
13 298 245 0 2 22
0 19 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
7100 0 0
2
44795.6 0
0
5 4081~
219 233 245 0 3 22
0 21 20 19
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndB
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3820 0 0
2
44795.6 0
0
5 4071~
219 143 209 0 3 22
0 23 22 21
0
0 0 624 0
4 4071
-7 -24 21 -16
3 OrB
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
7678 0 0
2
44795.6 0
0
14 Logic Display~
6 333 98 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90044e-315 0
0
9 Inverter~
13 285 113 0 2 22
0 25 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3178 0 0
2
5.90044e-315 0
0
5 4071~
219 209 113 0 3 22
0 27 26 25
0
0 0 624 0
4 4071
-7 -24 21 -16
3 Or1
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3409 0 0
2
5.90044e-315 0
0
5 4081~
219 149 72 0 3 22
0 29 28 27
0
0 0 624 0
4 4081
-7 -24 21 -16
4 And1
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3951 0 0
2
5.90044e-315 0
0
31
3 1 2 0 0 4224 0 16 15 0 0 4
414 563
445 563
445 568
458 568
3 1 3 0 0 4224 0 17 16 0 0 3
353 534
353 554
369 554
1 2 4 0 0 4224 0 1 16 0 0 4
54 602
356 602
356 572
369 572
2 1 5 0 0 4224 0 18 17 0 0 4
269 517
287 517
287 525
304 525
1 2 6 0 0 4224 0 2 17 0 0 4
53 564
277 564
277 543
304 543
3 1 7 0 0 4224 0 19 18 0 0 2
194 517
233 517
3 1 8 0 0 8320 0 20 19 0 0 4
134 483
140 483
140 508
149 508
1 2 9 0 0 4224 0 3 19 0 0 4
54 530
144 530
144 526
149 526
1 2 10 0 0 4224 0 4 20 0 0 4
54 497
74 497
74 492
88 492
1 1 11 0 0 4224 0 5 20 0 0 4
54 467
75 467
75 474
88 474
3 1 12 0 0 4224 0 24 21 0 0 4
297 374
319 374
319 379
327 379
4 2 13 0 0 4224 0 22 24 0 0 4
192 398
232 398
232 383
251 383
4 1 14 0 0 4224 0 23 24 0 0 4
182 344
227 344
227 365
251 365
1 3 15 0 0 4096 0 6 22 0 0 4
111 419
140 419
140 407
147 407
0 2 16 0 0 4096 0 0 22 18 0 3
122 372
122 398
147 398
0 1 17 0 0 4224 0 0 22 19 0 3
116 324
116 389
147 389
1 3 15 0 0 4224 0 6 23 0 0 3
111 419
111 353
131 353
1 2 16 0 0 8320 0 7 23 0 0 4
109 372
124 372
124 344
131 344
1 1 17 0 0 0 0 8 23 0 0 4
107 324
125 324
125 335
131 335
2 1 18 0 0 4224 0 26 25 0 0 4
319 245
340 245
340 249
351 249
3 1 19 0 0 4224 0 27 26 0 0 2
254 245
283 245
1 2 20 0 0 4224 0 9 27 0 0 4
107 284
195 284
195 254
209 254
3 1 21 0 0 8320 0 28 27 0 0 4
176 209
197 209
197 236
209 236
1 2 22 0 0 4224 0 10 28 0 0 4
106 234
124 234
124 218
130 218
1 1 23 0 0 4224 0 11 28 0 0 4
106 186
120 186
120 200
130 200
2 1 24 0 0 8320 0 30 29 0 0 3
306 113
306 116
333 116
3 1 25 0 0 4224 0 31 30 0 0 2
242 113
270 113
1 2 26 0 0 4224 0 12 31 0 0 3
99 128
196 128
196 122
3 1 27 0 0 4224 0 32 31 0 0 3
170 72
170 104
196 104
1 2 28 0 0 4224 0 14 32 0 0 4
100 91
117 91
117 81
125 81
1 1 29 0 0 4224 0 13 32 0 0 4
99 56
117 56
117 63
125 63
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
